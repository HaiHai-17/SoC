library verilog;
use verilog.vl_types.all;
entity system_nios2_qsys_0_nios2_performance_monitors is
end system_nios2_qsys_0_nios2_performance_monitors;
