library verilog;
use verilog.vl_types.all;
entity systemne_nios2_qsys_0_nios2_performance_monitors is
end systemne_nios2_qsys_0_nios2_performance_monitors;
