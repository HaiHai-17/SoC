library verilog;
use verilog.vl_types.all;
entity systemne_tb is
end systemne_tb;
