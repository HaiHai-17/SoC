library verilog;
use verilog.vl_types.all;
entity systemne is
    port(
        clk_clk         : in     vl_logic;
        reset_reset_n   : in     vl_logic
    );
end systemne;
