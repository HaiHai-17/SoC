library verilog;
use verilog.vl_types.all;
entity system_tb is
end system_tb;
