// nios_sys.v

// Generated using ACDS version 13.0sp1 232 at 2024.04.16.16:46:36

`timescale 1 ps / 1 ps
module nios_sys (
		input  wire        clk_clk,                             //                          clk.clk
		input  wire        reset_reset_n,                       //                        reset.reset_n
		output wire [6:0]  hex7_external_connection_export,     //     hex7_external_connection.export
		output wire [6:0]  hex6_external_connection_export,     //     hex6_external_connection.export
		output wire [6:0]  hex5_external_connection_export,     //     hex5_external_connection.export
		output wire [6:0]  hex4_external_connection_export,     //     hex4_external_connection.export
		output wire [6:0]  hex3_external_connection_export,     //     hex3_external_connection.export
		output wire [6:0]  hex2_external_connection_export,     //     hex2_external_connection.export
		output wire [6:0]  hex1_external_connection_export,     //     hex1_external_connection.export
		output wire [6:0]  hex0_external_connection_export,     //     hex0_external_connection.export
		output wire [17:0] ledr_external_connection_export,     //     ledr_external_connection.export
		input  wire [17:0] switch_external_connection_export,   //   switch_external_connection.export
		output wire [3:0]  ledg_external_connection_export,     //     ledg_external_connection.export
		input  wire [3:0]  key_external_connection_export,      //      key_external_connection.export
		output wire        lcd_rs_external_connection_export,   //   lcd_rs_external_connection.export
		output wire        lcd_rw_external_connection_export,   //   lcd_rw_external_connection.export
		output wire        lcd_en_external_connection_export,   //   lcd_en_external_connection.export
		output wire        lcd_blon_external_connection_export, // lcd_blon_external_connection.export
		output wire        lcd_on_external_connection_export,   //   lcd_on_external_connection.export
		output wire [7:0]  lcd_d_external_connection_export     //    lcd_d_external_connection.export
	);

	wire         nios2_qsys_0_instruction_master_waitrequest;                                                         // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                                                             // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                            // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                                                // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                  // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [16:0] nios2_qsys_0_data_master_address;                                                                    // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                      // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                       // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                   // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                 // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                           // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                  // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                        // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire  [12:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                          // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                       // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                            // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire         onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                            // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                         // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                       // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire   [1:0] switch_s1_translator_avalon_anti_slave_0_address;                                                    // switch_s1_translator:av_address -> switch:address
	wire  [31:0] switch_s1_translator_avalon_anti_slave_0_readdata;                                                   // switch:readdata -> switch_s1_translator:av_readdata
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_writedata;                                                    // ledr_s1_translator:av_writedata -> ledr:writedata
	wire   [1:0] ledr_s1_translator_avalon_anti_slave_0_address;                                                      // ledr_s1_translator:av_address -> ledr:address
	wire         ledr_s1_translator_avalon_anti_slave_0_chipselect;                                                   // ledr_s1_translator:av_chipselect -> ledr:chipselect
	wire         ledr_s1_translator_avalon_anti_slave_0_write;                                                        // ledr_s1_translator:av_write -> ledr:write_n
	wire  [31:0] ledr_s1_translator_avalon_anti_slave_0_readdata;                                                     // ledr:readdata -> ledr_s1_translator:av_readdata
	wire  [31:0] hex0_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex0_s1_translator:av_writedata -> hex0:writedata
	wire   [1:0] hex0_s1_translator_avalon_anti_slave_0_address;                                                      // hex0_s1_translator:av_address -> hex0:address
	wire         hex0_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex0_s1_translator:av_chipselect -> hex0:chipselect
	wire         hex0_s1_translator_avalon_anti_slave_0_write;                                                        // hex0_s1_translator:av_write -> hex0:write_n
	wire  [31:0] hex0_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex0:readdata -> hex0_s1_translator:av_readdata
	wire  [31:0] hex1_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex1_s1_translator:av_writedata -> hex1:writedata
	wire   [1:0] hex1_s1_translator_avalon_anti_slave_0_address;                                                      // hex1_s1_translator:av_address -> hex1:address
	wire         hex1_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex1_s1_translator:av_chipselect -> hex1:chipselect
	wire         hex1_s1_translator_avalon_anti_slave_0_write;                                                        // hex1_s1_translator:av_write -> hex1:write_n
	wire  [31:0] hex1_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex1:readdata -> hex1_s1_translator:av_readdata
	wire  [31:0] hex2_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex2_s1_translator:av_writedata -> hex2:writedata
	wire   [1:0] hex2_s1_translator_avalon_anti_slave_0_address;                                                      // hex2_s1_translator:av_address -> hex2:address
	wire         hex2_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex2_s1_translator:av_chipselect -> hex2:chipselect
	wire         hex2_s1_translator_avalon_anti_slave_0_write;                                                        // hex2_s1_translator:av_write -> hex2:write_n
	wire  [31:0] hex2_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex2:readdata -> hex2_s1_translator:av_readdata
	wire  [31:0] hex3_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex3_s1_translator:av_writedata -> hex3:writedata
	wire   [1:0] hex3_s1_translator_avalon_anti_slave_0_address;                                                      // hex3_s1_translator:av_address -> hex3:address
	wire         hex3_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex3_s1_translator:av_chipselect -> hex3:chipselect
	wire         hex3_s1_translator_avalon_anti_slave_0_write;                                                        // hex3_s1_translator:av_write -> hex3:write_n
	wire  [31:0] hex3_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex3:readdata -> hex3_s1_translator:av_readdata
	wire  [31:0] hex4_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex4_s1_translator:av_writedata -> hex4:writedata
	wire   [1:0] hex4_s1_translator_avalon_anti_slave_0_address;                                                      // hex4_s1_translator:av_address -> hex4:address
	wire         hex4_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex4_s1_translator:av_chipselect -> hex4:chipselect
	wire         hex4_s1_translator_avalon_anti_slave_0_write;                                                        // hex4_s1_translator:av_write -> hex4:write_n
	wire  [31:0] hex4_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex4:readdata -> hex4_s1_translator:av_readdata
	wire  [31:0] hex5_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex5_s1_translator:av_writedata -> hex5:writedata
	wire   [1:0] hex5_s1_translator_avalon_anti_slave_0_address;                                                      // hex5_s1_translator:av_address -> hex5:address
	wire         hex5_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex5_s1_translator:av_chipselect -> hex5:chipselect
	wire         hex5_s1_translator_avalon_anti_slave_0_write;                                                        // hex5_s1_translator:av_write -> hex5:write_n
	wire  [31:0] hex5_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex5:readdata -> hex5_s1_translator:av_readdata
	wire  [31:0] hex6_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex6_s1_translator:av_writedata -> hex6:writedata
	wire   [1:0] hex6_s1_translator_avalon_anti_slave_0_address;                                                      // hex6_s1_translator:av_address -> hex6:address
	wire         hex6_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex6_s1_translator:av_chipselect -> hex6:chipselect
	wire         hex6_s1_translator_avalon_anti_slave_0_write;                                                        // hex6_s1_translator:av_write -> hex6:write_n
	wire  [31:0] hex6_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex6:readdata -> hex6_s1_translator:av_readdata
	wire  [31:0] hex7_s1_translator_avalon_anti_slave_0_writedata;                                                    // hex7_s1_translator:av_writedata -> hex7:writedata
	wire   [1:0] hex7_s1_translator_avalon_anti_slave_0_address;                                                      // hex7_s1_translator:av_address -> hex7:address
	wire         hex7_s1_translator_avalon_anti_slave_0_chipselect;                                                   // hex7_s1_translator:av_chipselect -> hex7:chipselect
	wire         hex7_s1_translator_avalon_anti_slave_0_write;                                                        // hex7_s1_translator:av_write -> hex7:write_n
	wire  [31:0] hex7_s1_translator_avalon_anti_slave_0_readdata;                                                     // hex7:readdata -> hex7_s1_translator:av_readdata
	wire  [31:0] ledg_s1_translator_avalon_anti_slave_0_writedata;                                                    // ledg_s1_translator:av_writedata -> ledg:writedata
	wire   [1:0] ledg_s1_translator_avalon_anti_slave_0_address;                                                      // ledg_s1_translator:av_address -> ledg:address
	wire         ledg_s1_translator_avalon_anti_slave_0_chipselect;                                                   // ledg_s1_translator:av_chipselect -> ledg:chipselect
	wire         ledg_s1_translator_avalon_anti_slave_0_write;                                                        // ledg_s1_translator:av_write -> ledg:write_n
	wire  [31:0] ledg_s1_translator_avalon_anti_slave_0_readdata;                                                     // ledg:readdata -> ledg_s1_translator:av_readdata
	wire   [1:0] key_s1_translator_avalon_anti_slave_0_address;                                                       // key_s1_translator:av_address -> key:address
	wire  [31:0] key_s1_translator_avalon_anti_slave_0_readdata;                                                      // key:readdata -> key_s1_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                   // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                     // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire  [31:0] lcd_d_s1_translator_avalon_anti_slave_0_writedata;                                                   // lcd_d_s1_translator:av_writedata -> lcd_d:writedata
	wire   [1:0] lcd_d_s1_translator_avalon_anti_slave_0_address;                                                     // lcd_d_s1_translator:av_address -> lcd_d:address
	wire         lcd_d_s1_translator_avalon_anti_slave_0_chipselect;                                                  // lcd_d_s1_translator:av_chipselect -> lcd_d:chipselect
	wire         lcd_d_s1_translator_avalon_anti_slave_0_write;                                                       // lcd_d_s1_translator:av_write -> lcd_d:write_n
	wire  [31:0] lcd_d_s1_translator_avalon_anti_slave_0_readdata;                                                    // lcd_d:readdata -> lcd_d_s1_translator:av_readdata
	wire  [31:0] lcd_on_s1_translator_avalon_anti_slave_0_writedata;                                                  // lcd_on_s1_translator:av_writedata -> lcd_on:writedata
	wire   [1:0] lcd_on_s1_translator_avalon_anti_slave_0_address;                                                    // lcd_on_s1_translator:av_address -> lcd_on:address
	wire         lcd_on_s1_translator_avalon_anti_slave_0_chipselect;                                                 // lcd_on_s1_translator:av_chipselect -> lcd_on:chipselect
	wire         lcd_on_s1_translator_avalon_anti_slave_0_write;                                                      // lcd_on_s1_translator:av_write -> lcd_on:write_n
	wire  [31:0] lcd_on_s1_translator_avalon_anti_slave_0_readdata;                                                   // lcd_on:readdata -> lcd_on_s1_translator:av_readdata
	wire  [31:0] lcd_blon_s1_translator_avalon_anti_slave_0_writedata;                                                // lcd_blon_s1_translator:av_writedata -> lcd_blon:writedata
	wire   [1:0] lcd_blon_s1_translator_avalon_anti_slave_0_address;                                                  // lcd_blon_s1_translator:av_address -> lcd_blon:address
	wire         lcd_blon_s1_translator_avalon_anti_slave_0_chipselect;                                               // lcd_blon_s1_translator:av_chipselect -> lcd_blon:chipselect
	wire         lcd_blon_s1_translator_avalon_anti_slave_0_write;                                                    // lcd_blon_s1_translator:av_write -> lcd_blon:write_n
	wire  [31:0] lcd_blon_s1_translator_avalon_anti_slave_0_readdata;                                                 // lcd_blon:readdata -> lcd_blon_s1_translator:av_readdata
	wire  [31:0] lcd_en_s1_translator_avalon_anti_slave_0_writedata;                                                  // lcd_en_s1_translator:av_writedata -> lcd_en:writedata
	wire   [1:0] lcd_en_s1_translator_avalon_anti_slave_0_address;                                                    // lcd_en_s1_translator:av_address -> lcd_en:address
	wire         lcd_en_s1_translator_avalon_anti_slave_0_chipselect;                                                 // lcd_en_s1_translator:av_chipselect -> lcd_en:chipselect
	wire         lcd_en_s1_translator_avalon_anti_slave_0_write;                                                      // lcd_en_s1_translator:av_write -> lcd_en:write_n
	wire  [31:0] lcd_en_s1_translator_avalon_anti_slave_0_readdata;                                                   // lcd_en:readdata -> lcd_en_s1_translator:av_readdata
	wire  [31:0] lcd_rw_s1_translator_avalon_anti_slave_0_writedata;                                                  // lcd_rw_s1_translator:av_writedata -> lcd_rw:writedata
	wire   [1:0] lcd_rw_s1_translator_avalon_anti_slave_0_address;                                                    // lcd_rw_s1_translator:av_address -> lcd_rw:address
	wire         lcd_rw_s1_translator_avalon_anti_slave_0_chipselect;                                                 // lcd_rw_s1_translator:av_chipselect -> lcd_rw:chipselect
	wire         lcd_rw_s1_translator_avalon_anti_slave_0_write;                                                      // lcd_rw_s1_translator:av_write -> lcd_rw:write_n
	wire  [31:0] lcd_rw_s1_translator_avalon_anti_slave_0_readdata;                                                   // lcd_rw:readdata -> lcd_rw_s1_translator:av_readdata
	wire  [31:0] lcd_rs_s1_translator_avalon_anti_slave_0_writedata;                                                  // lcd_rs_s1_translator:av_writedata -> lcd_rs:writedata
	wire   [1:0] lcd_rs_s1_translator_avalon_anti_slave_0_address;                                                    // lcd_rs_s1_translator:av_address -> lcd_rs:address
	wire         lcd_rs_s1_translator_avalon_anti_slave_0_chipselect;                                                 // lcd_rs_s1_translator:av_chipselect -> lcd_rs:chipselect
	wire         lcd_rs_s1_translator_avalon_anti_slave_0_write;                                                      // lcd_rs_s1_translator:av_write -> lcd_rs:write_n
	wire  [31:0] lcd_rs_s1_translator_avalon_anti_slave_0_readdata;                                                   // lcd_rs:readdata -> lcd_rs_s1_translator:av_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [16:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [16:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [16:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [16:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire  [16:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire  [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                           // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // switch_s1_translator:uav_waitrequest -> switch_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // switch_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_s1_translator:uav_burstcount
	wire  [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // switch_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_s1_translator:uav_writedata
	wire  [16:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // switch_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_s1_translator:uav_address
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // switch_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_s1_translator:uav_write
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_s1_translator:uav_lock
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // switch_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_s1_translator:uav_read
	wire  [31:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // switch_s1_translator:uav_readdata -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // switch_s1_translator:uav_readdatavalid -> switch_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // switch_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_s1_translator:uav_debugaccess
	wire   [3:0] switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // switch_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_s1_translator:uav_byteenable
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // switch_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // ledr_s1_translator:uav_waitrequest -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledr_s1_translator:uav_burstcount
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // ledr_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledr_s1_translator:uav_writedata
	wire  [16:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // ledr_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledr_s1_translator:uav_address
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // ledr_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledr_s1_translator:uav_write
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledr_s1_translator:uav_lock
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledr_s1_translator:uav_read
	wire  [31:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // ledr_s1_translator:uav_readdata -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // ledr_s1_translator:uav_readdatavalid -> ledr_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledr_s1_translator:uav_debugaccess
	wire   [3:0] ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // ledr_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledr_s1_translator:uav_byteenable
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // ledr_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex0_s1_translator:uav_waitrequest -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex0_s1_translator:uav_burstcount
	wire  [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex0_s1_translator:uav_writedata
	wire  [16:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex0_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex0_s1_translator:uav_address
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex0_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex0_s1_translator:uav_write
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex0_s1_translator:uav_lock
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex0_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex0_s1_translator:uav_read
	wire  [31:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex0_s1_translator:uav_readdata -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex0_s1_translator:uav_readdatavalid -> hex0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex0_s1_translator:uav_debugaccess
	wire   [3:0] hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex0_s1_translator:uav_byteenable
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex1_s1_translator:uav_waitrequest -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex1_s1_translator:uav_burstcount
	wire  [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex1_s1_translator:uav_writedata
	wire  [16:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex1_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex1_s1_translator:uav_address
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex1_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex1_s1_translator:uav_write
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex1_s1_translator:uav_lock
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex1_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex1_s1_translator:uav_read
	wire  [31:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex1_s1_translator:uav_readdata -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex1_s1_translator:uav_readdatavalid -> hex1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex1_s1_translator:uav_debugaccess
	wire   [3:0] hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex1_s1_translator:uav_byteenable
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex2_s1_translator:uav_waitrequest -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex2_s1_translator:uav_burstcount
	wire  [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex2_s1_translator:uav_writedata
	wire  [16:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex2_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex2_s1_translator:uav_address
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex2_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex2_s1_translator:uav_write
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex2_s1_translator:uav_lock
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex2_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex2_s1_translator:uav_read
	wire  [31:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex2_s1_translator:uav_readdata -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex2_s1_translator:uav_readdatavalid -> hex2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex2_s1_translator:uav_debugaccess
	wire   [3:0] hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex2_s1_translator:uav_byteenable
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex3_s1_translator:uav_waitrequest -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex3_s1_translator:uav_burstcount
	wire  [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex3_s1_translator:uav_writedata
	wire  [16:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex3_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex3_s1_translator:uav_address
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex3_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex3_s1_translator:uav_write
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex3_s1_translator:uav_lock
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex3_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex3_s1_translator:uav_read
	wire  [31:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex3_s1_translator:uav_readdata -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex3_s1_translator:uav_readdatavalid -> hex3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex3_s1_translator:uav_debugaccess
	wire   [3:0] hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex3_s1_translator:uav_byteenable
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex4_s1_translator:uav_waitrequest -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex4_s1_translator:uav_burstcount
	wire  [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex4_s1_translator:uav_writedata
	wire  [16:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex4_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex4_s1_translator:uav_address
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex4_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex4_s1_translator:uav_write
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex4_s1_translator:uav_lock
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex4_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex4_s1_translator:uav_read
	wire  [31:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex4_s1_translator:uav_readdata -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex4_s1_translator:uav_readdatavalid -> hex4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex4_s1_translator:uav_debugaccess
	wire   [3:0] hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex4_s1_translator:uav_byteenable
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex5_s1_translator:uav_waitrequest -> hex5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex5_s1_translator:uav_burstcount
	wire  [31:0] hex5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex5_s1_translator:uav_writedata
	wire  [16:0] hex5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex5_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex5_s1_translator:uav_address
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex5_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex5_s1_translator:uav_write
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex5_s1_translator:uav_lock
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex5_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex5_s1_translator:uav_read
	wire  [31:0] hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex5_s1_translator:uav_readdata -> hex5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex5_s1_translator:uav_readdatavalid -> hex5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex5_s1_translator:uav_debugaccess
	wire   [3:0] hex5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex5_s1_translator:uav_byteenable
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex6_s1_translator:uav_waitrequest -> hex6_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex6_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex6_s1_translator:uav_burstcount
	wire  [31:0] hex6_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex6_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex6_s1_translator:uav_writedata
	wire  [16:0] hex6_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex6_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex6_s1_translator:uav_address
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex6_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex6_s1_translator:uav_write
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex6_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex6_s1_translator:uav_lock
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex6_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex6_s1_translator:uav_read
	wire  [31:0] hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex6_s1_translator:uav_readdata -> hex6_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex6_s1_translator:uav_readdatavalid -> hex6_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex6_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex6_s1_translator:uav_debugaccess
	wire   [3:0] hex6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex6_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex6_s1_translator:uav_byteenable
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex6_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex6_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex6_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex6_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex6_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex6_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex6_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex6_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // hex7_s1_translator:uav_waitrequest -> hex7_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] hex7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // hex7_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hex7_s1_translator:uav_burstcount
	wire  [31:0] hex7_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // hex7_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hex7_s1_translator:uav_writedata
	wire  [16:0] hex7_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // hex7_s1_translator_avalon_universal_slave_0_agent:m0_address -> hex7_s1_translator:uav_address
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // hex7_s1_translator_avalon_universal_slave_0_agent:m0_write -> hex7_s1_translator:uav_write
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // hex7_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hex7_s1_translator:uav_lock
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // hex7_s1_translator_avalon_universal_slave_0_agent:m0_read -> hex7_s1_translator:uav_read
	wire  [31:0] hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // hex7_s1_translator:uav_readdata -> hex7_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // hex7_s1_translator:uav_readdatavalid -> hex7_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // hex7_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hex7_s1_translator:uav_debugaccess
	wire   [3:0] hex7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // hex7_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hex7_s1_translator:uav_byteenable
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // hex7_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // hex7_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // hex7_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // hex7_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hex7_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hex7_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hex7_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // hex7_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hex7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // ledg_s1_translator:uav_waitrequest -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // ledg_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ledg_s1_translator:uav_burstcount
	wire  [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // ledg_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ledg_s1_translator:uav_writedata
	wire  [16:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // ledg_s1_translator_avalon_universal_slave_0_agent:m0_address -> ledg_s1_translator:uav_address
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // ledg_s1_translator_avalon_universal_slave_0_agent:m0_write -> ledg_s1_translator:uav_write
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // ledg_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ledg_s1_translator:uav_lock
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // ledg_s1_translator_avalon_universal_slave_0_agent:m0_read -> ledg_s1_translator:uav_read
	wire  [31:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // ledg_s1_translator:uav_readdata -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // ledg_s1_translator:uav_readdatavalid -> ledg_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // ledg_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ledg_s1_translator:uav_debugaccess
	wire   [3:0] ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // ledg_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ledg_s1_translator:uav_byteenable
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // ledg_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // key_s1_translator:uav_waitrequest -> key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> key_s1_translator:uav_burstcount
	wire  [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> key_s1_translator:uav_writedata
	wire  [16:0] key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // key_s1_translator_avalon_universal_slave_0_agent:m0_address -> key_s1_translator:uav_address
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // key_s1_translator_avalon_universal_slave_0_agent:m0_write -> key_s1_translator:uav_write
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> key_s1_translator:uav_lock
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // key_s1_translator_avalon_universal_slave_0_agent:m0_read -> key_s1_translator:uav_read
	wire  [31:0] key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // key_s1_translator:uav_readdata -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // key_s1_translator:uav_readdatavalid -> key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> key_s1_translator:uav_debugaccess
	wire   [3:0] key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> key_s1_translator:uav_byteenable
	wire         key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [16:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // lcd_d_s1_translator:uav_waitrequest -> lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_d_s1_translator:uav_burstcount
	wire  [31:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_d_s1_translator:uav_writedata
	wire  [16:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_d_s1_translator:uav_address
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_d_s1_translator:uav_write
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_d_s1_translator:uav_lock
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_d_s1_translator:uav_read
	wire  [31:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // lcd_d_s1_translator:uav_readdata -> lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // lcd_d_s1_translator:uav_readdatavalid -> lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_d_s1_translator:uav_debugaccess
	wire   [3:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // lcd_d_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_d_s1_translator:uav_byteenable
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // lcd_d_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // lcd_on_s1_translator:uav_waitrequest -> lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_on_s1_translator:uav_burstcount
	wire  [31:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_on_s1_translator:uav_writedata
	wire  [16:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_on_s1_translator:uav_address
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_on_s1_translator:uav_write
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_on_s1_translator:uav_lock
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_on_s1_translator:uav_read
	wire  [31:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // lcd_on_s1_translator:uav_readdata -> lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // lcd_on_s1_translator:uav_readdatavalid -> lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_on_s1_translator:uav_debugaccess
	wire   [3:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // lcd_on_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_on_s1_translator:uav_byteenable
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // lcd_on_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // lcd_blon_s1_translator:uav_waitrequest -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_blon_s1_translator:uav_burstcount
	wire  [31:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_blon_s1_translator:uav_writedata
	wire  [16:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_blon_s1_translator:uav_address
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_blon_s1_translator:uav_write
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_blon_s1_translator:uav_lock
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_blon_s1_translator:uav_read
	wire  [31:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // lcd_blon_s1_translator:uav_readdata -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // lcd_blon_s1_translator:uav_readdatavalid -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_blon_s1_translator:uav_debugaccess
	wire   [3:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // lcd_blon_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_blon_s1_translator:uav_byteenable
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // lcd_en_s1_translator:uav_waitrequest -> lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_en_s1_translator:uav_burstcount
	wire  [31:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_en_s1_translator:uav_writedata
	wire  [16:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_en_s1_translator:uav_address
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_en_s1_translator:uav_write
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_en_s1_translator:uav_lock
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_en_s1_translator:uav_read
	wire  [31:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // lcd_en_s1_translator:uav_readdata -> lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // lcd_en_s1_translator:uav_readdatavalid -> lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_en_s1_translator:uav_debugaccess
	wire   [3:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // lcd_en_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_en_s1_translator:uav_byteenable
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // lcd_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // lcd_rw_s1_translator:uav_waitrequest -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_rw_s1_translator:uav_burstcount
	wire  [31:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_rw_s1_translator:uav_writedata
	wire  [16:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_rw_s1_translator:uav_address
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_rw_s1_translator:uav_write
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_rw_s1_translator:uav_lock
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_rw_s1_translator:uav_read
	wire  [31:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // lcd_rw_s1_translator:uav_readdata -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // lcd_rw_s1_translator:uav_readdatavalid -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_rw_s1_translator:uav_debugaccess
	wire   [3:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // lcd_rw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_rw_s1_translator:uav_byteenable
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // lcd_rs_s1_translator:uav_waitrequest -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_rs_s1_translator:uav_burstcount
	wire  [31:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_rs_s1_translator:uav_writedata
	wire  [16:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_rs_s1_translator:uav_address
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_rs_s1_translator:uav_write
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_rs_s1_translator:uav_lock
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_rs_s1_translator:uav_read
	wire  [31:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // lcd_rs_s1_translator:uav_readdata -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // lcd_rs_s1_translator:uav_readdatavalid -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_rs_s1_translator:uav_debugaccess
	wire   [3:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // lcd_rs_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_rs_s1_translator:uav_byteenable
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [94:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [94:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [93:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [93:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [93:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [93:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_001:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [93:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_002:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // switch_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // switch_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // switch_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [93:0] switch_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // switch_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         switch_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_003:sink_ready -> switch_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // ledr_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // ledr_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // ledr_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [93:0] ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // ledr_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_004:sink_ready -> ledr_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [93:0] hex0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_005:sink_ready -> hex0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [93:0] hex1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_006:sink_ready -> hex1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [93:0] hex2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_007:sink_ready -> hex2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [93:0] hex3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_008:sink_ready -> hex3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [93:0] hex4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_009:sink_ready -> hex4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [93:0] hex5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         hex5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_010:sink_ready -> hex5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex6_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex6_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex6_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [93:0] hex6_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex6_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         hex6_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_011:sink_ready -> hex6_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // hex7_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // hex7_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // hex7_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [93:0] hex7_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // hex7_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         hex7_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_012:sink_ready -> hex7_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // ledg_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // ledg_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // ledg_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [93:0] ledg_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // ledg_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_013:sink_ready -> ledg_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire         key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire         key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [93:0] key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire         key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_014:sink_ready -> key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [93:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_015:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // lcd_d_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // lcd_d_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // lcd_d_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [93:0] lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // lcd_d_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire         lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_016:sink_ready -> lcd_d_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // lcd_on_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // lcd_on_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // lcd_on_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [93:0] lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // lcd_on_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire         lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_017:sink_ready -> lcd_on_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [93:0] lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // lcd_blon_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire         lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_018:sink_ready -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // lcd_en_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // lcd_en_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // lcd_en_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire  [93:0] lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // lcd_en_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire         lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_019:sink_ready -> lcd_en_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [93:0] lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // lcd_rw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire         lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_020:sink_ready -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	wire  [93:0] lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // lcd_rs_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	wire         lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_021:sink_ready -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, cmd_xbar_mux_015:reset, cmd_xbar_mux_016:reset, cmd_xbar_mux_017:reset, cmd_xbar_mux_018:reset, cmd_xbar_mux_019:reset, cmd_xbar_mux_020:reset, cmd_xbar_mux_021:reset, hex0:reset_n, hex0_s1_translator:reset, hex0_s1_translator_avalon_universal_slave_0_agent:reset, hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex1:reset_n, hex1_s1_translator:reset, hex1_s1_translator_avalon_universal_slave_0_agent:reset, hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex2:reset_n, hex2_s1_translator:reset, hex2_s1_translator_avalon_universal_slave_0_agent:reset, hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex3:reset_n, hex3_s1_translator:reset, hex3_s1_translator_avalon_universal_slave_0_agent:reset, hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex4:reset_n, hex4_s1_translator:reset, hex4_s1_translator_avalon_universal_slave_0_agent:reset, hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex5:reset_n, hex5_s1_translator:reset, hex5_s1_translator_avalon_universal_slave_0_agent:reset, hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex6:reset_n, hex6_s1_translator:reset, hex6_s1_translator_avalon_universal_slave_0_agent:reset, hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hex7:reset_n, hex7_s1_translator:reset, hex7_s1_translator_avalon_universal_slave_0_agent:reset, hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, key:reset_n, key_s1_translator:reset, key_s1_translator_avalon_universal_slave_0_agent:reset, key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_blon:reset_n, lcd_blon_s1_translator:reset, lcd_blon_s1_translator_avalon_universal_slave_0_agent:reset, lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_d:reset_n, lcd_d_s1_translator:reset, lcd_d_s1_translator_avalon_universal_slave_0_agent:reset, lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_en:reset_n, lcd_en_s1_translator:reset, lcd_en_s1_translator_avalon_universal_slave_0_agent:reset, lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_on:reset_n, lcd_on_s1_translator:reset, lcd_on_s1_translator_avalon_universal_slave_0_agent:reset, lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_rs:reset_n, lcd_rs_s1_translator:reset, lcd_rs_s1_translator_avalon_universal_slave_0_agent:reset, lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_rw:reset_n, lcd_rw_s1_translator:reset, lcd_rw_s1_translator_avalon_universal_slave_0_agent:reset, lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledg:reset_n, ledg_s1_translator:reset, ledg_s1_translator_avalon_universal_slave_0_agent:reset, ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ledr:reset_n, ledr_s1_translator:reset, ledr_s1_translator_avalon_universal_slave_0_agent:reset, ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, switch:reset_n, switch_s1_translator:reset, switch_s1_translator_avalon_universal_slave_0_agent:reset, switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_reset_out_reset_req;                                                                  // rst_controller:reset_req -> onchip_memory2_0:reset_req
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                          // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [21:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [21:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire  [21:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_src3_endofpacket;                                                                     // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                           // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                   // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src3_data;                                                                            // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire  [21:0] cmd_xbar_demux_src3_channel;                                                                         // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire         cmd_xbar_demux_src3_ready;                                                                           // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire         cmd_xbar_demux_src4_endofpacket;                                                                     // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                           // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                   // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src4_data;                                                                            // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire  [21:0] cmd_xbar_demux_src4_channel;                                                                         // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire         cmd_xbar_demux_src4_ready;                                                                           // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire         cmd_xbar_demux_src5_endofpacket;                                                                     // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire         cmd_xbar_demux_src5_valid;                                                                           // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire         cmd_xbar_demux_src5_startofpacket;                                                                   // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src5_data;                                                                            // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire  [21:0] cmd_xbar_demux_src5_channel;                                                                         // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire         cmd_xbar_demux_src5_ready;                                                                           // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire         cmd_xbar_demux_src6_endofpacket;                                                                     // cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire         cmd_xbar_demux_src6_valid;                                                                           // cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	wire         cmd_xbar_demux_src6_startofpacket;                                                                   // cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src6_data;                                                                            // cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	wire  [21:0] cmd_xbar_demux_src6_channel;                                                                         // cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	wire         cmd_xbar_demux_src6_ready;                                                                           // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	wire         cmd_xbar_demux_src7_endofpacket;                                                                     // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire         cmd_xbar_demux_src7_valid;                                                                           // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire         cmd_xbar_demux_src7_startofpacket;                                                                   // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src7_data;                                                                            // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire  [21:0] cmd_xbar_demux_src7_channel;                                                                         // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire         cmd_xbar_demux_src7_ready;                                                                           // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire         cmd_xbar_demux_src8_endofpacket;                                                                     // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire         cmd_xbar_demux_src8_valid;                                                                           // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire         cmd_xbar_demux_src8_startofpacket;                                                                   // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src8_data;                                                                            // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire  [21:0] cmd_xbar_demux_src8_channel;                                                                         // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire         cmd_xbar_demux_src8_ready;                                                                           // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire         cmd_xbar_demux_src9_endofpacket;                                                                     // cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire         cmd_xbar_demux_src9_valid;                                                                           // cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire         cmd_xbar_demux_src9_startofpacket;                                                                   // cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src9_data;                                                                            // cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	wire  [21:0] cmd_xbar_demux_src9_channel;                                                                         // cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire         cmd_xbar_demux_src9_ready;                                                                           // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire         cmd_xbar_demux_src10_endofpacket;                                                                    // cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire         cmd_xbar_demux_src10_valid;                                                                          // cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire         cmd_xbar_demux_src10_startofpacket;                                                                  // cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src10_data;                                                                           // cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	wire  [21:0] cmd_xbar_demux_src10_channel;                                                                        // cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire         cmd_xbar_demux_src10_ready;                                                                          // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire         cmd_xbar_demux_src11_endofpacket;                                                                    // cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	wire         cmd_xbar_demux_src11_valid;                                                                          // cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	wire         cmd_xbar_demux_src11_startofpacket;                                                                  // cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src11_data;                                                                           // cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	wire  [21:0] cmd_xbar_demux_src11_channel;                                                                        // cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	wire         cmd_xbar_demux_src11_ready;                                                                          // cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	wire         cmd_xbar_demux_src12_endofpacket;                                                                    // cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire         cmd_xbar_demux_src12_valid;                                                                          // cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	wire         cmd_xbar_demux_src12_startofpacket;                                                                  // cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src12_data;                                                                           // cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	wire  [21:0] cmd_xbar_demux_src12_channel;                                                                        // cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	wire         cmd_xbar_demux_src12_ready;                                                                          // cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	wire         cmd_xbar_demux_src13_endofpacket;                                                                    // cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire         cmd_xbar_demux_src13_valid;                                                                          // cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire         cmd_xbar_demux_src13_startofpacket;                                                                  // cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src13_data;                                                                           // cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	wire  [21:0] cmd_xbar_demux_src13_channel;                                                                        // cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire         cmd_xbar_demux_src13_ready;                                                                          // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	wire         cmd_xbar_demux_src14_endofpacket;                                                                    // cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	wire         cmd_xbar_demux_src14_valid;                                                                          // cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	wire         cmd_xbar_demux_src14_startofpacket;                                                                  // cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src14_data;                                                                           // cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	wire  [21:0] cmd_xbar_demux_src14_channel;                                                                        // cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	wire         cmd_xbar_demux_src14_ready;                                                                          // cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	wire         cmd_xbar_demux_src15_endofpacket;                                                                    // cmd_xbar_demux:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire         cmd_xbar_demux_src15_valid;                                                                          // cmd_xbar_demux:src15_valid -> cmd_xbar_mux_015:sink0_valid
	wire         cmd_xbar_demux_src15_startofpacket;                                                                  // cmd_xbar_demux:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src15_data;                                                                           // cmd_xbar_demux:src15_data -> cmd_xbar_mux_015:sink0_data
	wire  [21:0] cmd_xbar_demux_src15_channel;                                                                        // cmd_xbar_demux:src15_channel -> cmd_xbar_mux_015:sink0_channel
	wire         cmd_xbar_demux_src15_ready;                                                                          // cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux:src15_ready
	wire         cmd_xbar_demux_src16_endofpacket;                                                                    // cmd_xbar_demux:src16_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	wire         cmd_xbar_demux_src16_valid;                                                                          // cmd_xbar_demux:src16_valid -> cmd_xbar_mux_016:sink0_valid
	wire         cmd_xbar_demux_src16_startofpacket;                                                                  // cmd_xbar_demux:src16_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src16_data;                                                                           // cmd_xbar_demux:src16_data -> cmd_xbar_mux_016:sink0_data
	wire  [21:0] cmd_xbar_demux_src16_channel;                                                                        // cmd_xbar_demux:src16_channel -> cmd_xbar_mux_016:sink0_channel
	wire         cmd_xbar_demux_src16_ready;                                                                          // cmd_xbar_mux_016:sink0_ready -> cmd_xbar_demux:src16_ready
	wire         cmd_xbar_demux_src17_endofpacket;                                                                    // cmd_xbar_demux:src17_endofpacket -> cmd_xbar_mux_017:sink0_endofpacket
	wire         cmd_xbar_demux_src17_valid;                                                                          // cmd_xbar_demux:src17_valid -> cmd_xbar_mux_017:sink0_valid
	wire         cmd_xbar_demux_src17_startofpacket;                                                                  // cmd_xbar_demux:src17_startofpacket -> cmd_xbar_mux_017:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src17_data;                                                                           // cmd_xbar_demux:src17_data -> cmd_xbar_mux_017:sink0_data
	wire  [21:0] cmd_xbar_demux_src17_channel;                                                                        // cmd_xbar_demux:src17_channel -> cmd_xbar_mux_017:sink0_channel
	wire         cmd_xbar_demux_src17_ready;                                                                          // cmd_xbar_mux_017:sink0_ready -> cmd_xbar_demux:src17_ready
	wire         cmd_xbar_demux_src18_endofpacket;                                                                    // cmd_xbar_demux:src18_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	wire         cmd_xbar_demux_src18_valid;                                                                          // cmd_xbar_demux:src18_valid -> cmd_xbar_mux_018:sink0_valid
	wire         cmd_xbar_demux_src18_startofpacket;                                                                  // cmd_xbar_demux:src18_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src18_data;                                                                           // cmd_xbar_demux:src18_data -> cmd_xbar_mux_018:sink0_data
	wire  [21:0] cmd_xbar_demux_src18_channel;                                                                        // cmd_xbar_demux:src18_channel -> cmd_xbar_mux_018:sink0_channel
	wire         cmd_xbar_demux_src18_ready;                                                                          // cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux:src18_ready
	wire         cmd_xbar_demux_src19_endofpacket;                                                                    // cmd_xbar_demux:src19_endofpacket -> cmd_xbar_mux_019:sink0_endofpacket
	wire         cmd_xbar_demux_src19_valid;                                                                          // cmd_xbar_demux:src19_valid -> cmd_xbar_mux_019:sink0_valid
	wire         cmd_xbar_demux_src19_startofpacket;                                                                  // cmd_xbar_demux:src19_startofpacket -> cmd_xbar_mux_019:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src19_data;                                                                           // cmd_xbar_demux:src19_data -> cmd_xbar_mux_019:sink0_data
	wire  [21:0] cmd_xbar_demux_src19_channel;                                                                        // cmd_xbar_demux:src19_channel -> cmd_xbar_mux_019:sink0_channel
	wire         cmd_xbar_demux_src19_ready;                                                                          // cmd_xbar_mux_019:sink0_ready -> cmd_xbar_demux:src19_ready
	wire         cmd_xbar_demux_src20_endofpacket;                                                                    // cmd_xbar_demux:src20_endofpacket -> cmd_xbar_mux_020:sink0_endofpacket
	wire         cmd_xbar_demux_src20_valid;                                                                          // cmd_xbar_demux:src20_valid -> cmd_xbar_mux_020:sink0_valid
	wire         cmd_xbar_demux_src20_startofpacket;                                                                  // cmd_xbar_demux:src20_startofpacket -> cmd_xbar_mux_020:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src20_data;                                                                           // cmd_xbar_demux:src20_data -> cmd_xbar_mux_020:sink0_data
	wire  [21:0] cmd_xbar_demux_src20_channel;                                                                        // cmd_xbar_demux:src20_channel -> cmd_xbar_mux_020:sink0_channel
	wire         cmd_xbar_demux_src20_ready;                                                                          // cmd_xbar_mux_020:sink0_ready -> cmd_xbar_demux:src20_ready
	wire         cmd_xbar_demux_src21_endofpacket;                                                                    // cmd_xbar_demux:src21_endofpacket -> cmd_xbar_mux_021:sink0_endofpacket
	wire         cmd_xbar_demux_src21_valid;                                                                          // cmd_xbar_demux:src21_valid -> cmd_xbar_mux_021:sink0_valid
	wire         cmd_xbar_demux_src21_startofpacket;                                                                  // cmd_xbar_demux:src21_startofpacket -> cmd_xbar_mux_021:sink0_startofpacket
	wire  [93:0] cmd_xbar_demux_src21_data;                                                                           // cmd_xbar_demux:src21_data -> cmd_xbar_mux_021:sink0_data
	wire  [21:0] cmd_xbar_demux_src21_channel;                                                                        // cmd_xbar_demux:src21_channel -> cmd_xbar_mux_021:sink0_channel
	wire         cmd_xbar_demux_src21_ready;                                                                          // cmd_xbar_mux_021:sink0_ready -> cmd_xbar_demux:src21_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire         cmd_xbar_demux_001_src3_ready;                                                                       // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire         cmd_xbar_demux_001_src4_ready;                                                                       // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire         cmd_xbar_demux_001_src5_ready;                                                                       // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	wire         cmd_xbar_demux_001_src6_ready;                                                                       // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire         cmd_xbar_demux_001_src7_ready;                                                                       // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                                 // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                       // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                               // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src8_data;                                                                        // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src8_channel;                                                                     // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	wire         cmd_xbar_demux_001_src8_ready;                                                                       // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                                 // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                       // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                               // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src9_data;                                                                        // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src9_channel;                                                                     // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	wire         cmd_xbar_demux_001_src9_ready;                                                                       // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                                // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                      // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                              // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src10_data;                                                                       // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src10_channel;                                                                    // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	wire         cmd_xbar_demux_001_src10_ready;                                                                      // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                                // cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                      // cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink1_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                              // cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src11_data;                                                                       // cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src11_channel;                                                                    // cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink1_channel
	wire         cmd_xbar_demux_001_src11_ready;                                                                      // cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_001:src11_ready
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                                // cmd_xbar_demux_001:src12_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                      // cmd_xbar_demux_001:src12_valid -> cmd_xbar_mux_012:sink1_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                              // cmd_xbar_demux_001:src12_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src12_data;                                                                       // cmd_xbar_demux_001:src12_data -> cmd_xbar_mux_012:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src12_channel;                                                                    // cmd_xbar_demux_001:src12_channel -> cmd_xbar_mux_012:sink1_channel
	wire         cmd_xbar_demux_001_src12_ready;                                                                      // cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_001:src12_ready
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                                // cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                      // cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink1_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                              // cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src13_data;                                                                       // cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src13_channel;                                                                    // cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink1_channel
	wire         cmd_xbar_demux_001_src13_ready;                                                                      // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src13_ready
	wire         cmd_xbar_demux_001_src14_endofpacket;                                                                // cmd_xbar_demux_001:src14_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	wire         cmd_xbar_demux_001_src14_valid;                                                                      // cmd_xbar_demux_001:src14_valid -> cmd_xbar_mux_014:sink1_valid
	wire         cmd_xbar_demux_001_src14_startofpacket;                                                              // cmd_xbar_demux_001:src14_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src14_data;                                                                       // cmd_xbar_demux_001:src14_data -> cmd_xbar_mux_014:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src14_channel;                                                                    // cmd_xbar_demux_001:src14_channel -> cmd_xbar_mux_014:sink1_channel
	wire         cmd_xbar_demux_001_src14_ready;                                                                      // cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_001:src14_ready
	wire         cmd_xbar_demux_001_src15_endofpacket;                                                                // cmd_xbar_demux_001:src15_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire         cmd_xbar_demux_001_src15_valid;                                                                      // cmd_xbar_demux_001:src15_valid -> cmd_xbar_mux_015:sink1_valid
	wire         cmd_xbar_demux_001_src15_startofpacket;                                                              // cmd_xbar_demux_001:src15_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src15_data;                                                                       // cmd_xbar_demux_001:src15_data -> cmd_xbar_mux_015:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src15_channel;                                                                    // cmd_xbar_demux_001:src15_channel -> cmd_xbar_mux_015:sink1_channel
	wire         cmd_xbar_demux_001_src15_ready;                                                                      // cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_001:src15_ready
	wire         cmd_xbar_demux_001_src16_endofpacket;                                                                // cmd_xbar_demux_001:src16_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	wire         cmd_xbar_demux_001_src16_valid;                                                                      // cmd_xbar_demux_001:src16_valid -> cmd_xbar_mux_016:sink1_valid
	wire         cmd_xbar_demux_001_src16_startofpacket;                                                              // cmd_xbar_demux_001:src16_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src16_data;                                                                       // cmd_xbar_demux_001:src16_data -> cmd_xbar_mux_016:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src16_channel;                                                                    // cmd_xbar_demux_001:src16_channel -> cmd_xbar_mux_016:sink1_channel
	wire         cmd_xbar_demux_001_src16_ready;                                                                      // cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_001:src16_ready
	wire         cmd_xbar_demux_001_src17_endofpacket;                                                                // cmd_xbar_demux_001:src17_endofpacket -> cmd_xbar_mux_017:sink1_endofpacket
	wire         cmd_xbar_demux_001_src17_valid;                                                                      // cmd_xbar_demux_001:src17_valid -> cmd_xbar_mux_017:sink1_valid
	wire         cmd_xbar_demux_001_src17_startofpacket;                                                              // cmd_xbar_demux_001:src17_startofpacket -> cmd_xbar_mux_017:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src17_data;                                                                       // cmd_xbar_demux_001:src17_data -> cmd_xbar_mux_017:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src17_channel;                                                                    // cmd_xbar_demux_001:src17_channel -> cmd_xbar_mux_017:sink1_channel
	wire         cmd_xbar_demux_001_src17_ready;                                                                      // cmd_xbar_mux_017:sink1_ready -> cmd_xbar_demux_001:src17_ready
	wire         cmd_xbar_demux_001_src18_endofpacket;                                                                // cmd_xbar_demux_001:src18_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	wire         cmd_xbar_demux_001_src18_valid;                                                                      // cmd_xbar_demux_001:src18_valid -> cmd_xbar_mux_018:sink1_valid
	wire         cmd_xbar_demux_001_src18_startofpacket;                                                              // cmd_xbar_demux_001:src18_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src18_data;                                                                       // cmd_xbar_demux_001:src18_data -> cmd_xbar_mux_018:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src18_channel;                                                                    // cmd_xbar_demux_001:src18_channel -> cmd_xbar_mux_018:sink1_channel
	wire         cmd_xbar_demux_001_src18_ready;                                                                      // cmd_xbar_mux_018:sink1_ready -> cmd_xbar_demux_001:src18_ready
	wire         cmd_xbar_demux_001_src19_endofpacket;                                                                // cmd_xbar_demux_001:src19_endofpacket -> cmd_xbar_mux_019:sink1_endofpacket
	wire         cmd_xbar_demux_001_src19_valid;                                                                      // cmd_xbar_demux_001:src19_valid -> cmd_xbar_mux_019:sink1_valid
	wire         cmd_xbar_demux_001_src19_startofpacket;                                                              // cmd_xbar_demux_001:src19_startofpacket -> cmd_xbar_mux_019:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src19_data;                                                                       // cmd_xbar_demux_001:src19_data -> cmd_xbar_mux_019:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src19_channel;                                                                    // cmd_xbar_demux_001:src19_channel -> cmd_xbar_mux_019:sink1_channel
	wire         cmd_xbar_demux_001_src19_ready;                                                                      // cmd_xbar_mux_019:sink1_ready -> cmd_xbar_demux_001:src19_ready
	wire         cmd_xbar_demux_001_src20_endofpacket;                                                                // cmd_xbar_demux_001:src20_endofpacket -> cmd_xbar_mux_020:sink1_endofpacket
	wire         cmd_xbar_demux_001_src20_valid;                                                                      // cmd_xbar_demux_001:src20_valid -> cmd_xbar_mux_020:sink1_valid
	wire         cmd_xbar_demux_001_src20_startofpacket;                                                              // cmd_xbar_demux_001:src20_startofpacket -> cmd_xbar_mux_020:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src20_data;                                                                       // cmd_xbar_demux_001:src20_data -> cmd_xbar_mux_020:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src20_channel;                                                                    // cmd_xbar_demux_001:src20_channel -> cmd_xbar_mux_020:sink1_channel
	wire         cmd_xbar_demux_001_src20_ready;                                                                      // cmd_xbar_mux_020:sink1_ready -> cmd_xbar_demux_001:src20_ready
	wire         cmd_xbar_demux_001_src21_endofpacket;                                                                // cmd_xbar_demux_001:src21_endofpacket -> cmd_xbar_mux_021:sink1_endofpacket
	wire         cmd_xbar_demux_001_src21_valid;                                                                      // cmd_xbar_demux_001:src21_valid -> cmd_xbar_mux_021:sink1_valid
	wire         cmd_xbar_demux_001_src21_startofpacket;                                                              // cmd_xbar_demux_001:src21_startofpacket -> cmd_xbar_mux_021:sink1_startofpacket
	wire  [93:0] cmd_xbar_demux_001_src21_data;                                                                       // cmd_xbar_demux_001:src21_data -> cmd_xbar_mux_021:sink1_data
	wire  [21:0] cmd_xbar_demux_001_src21_channel;                                                                    // cmd_xbar_demux_001:src21_channel -> cmd_xbar_mux_021:sink1_channel
	wire         cmd_xbar_demux_001_src21_ready;                                                                      // cmd_xbar_mux_021:sink1_ready -> cmd_xbar_demux_001:src21_ready
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [21:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [93:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [21:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [21:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [93:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [21:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [93:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire  [21:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [93:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire  [21:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [93:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire  [21:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_003_src1_endofpacket;                                                                 // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src1_valid;                                                                       // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src1_startofpacket;                                                               // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [93:0] rsp_xbar_demux_003_src1_data;                                                                        // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire  [21:0] rsp_xbar_demux_003_src1_channel;                                                                     // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src1_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [93:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire  [21:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_004_src1_endofpacket;                                                                 // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src1_valid;                                                                       // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src1_startofpacket;                                                               // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [93:0] rsp_xbar_demux_004_src1_data;                                                                        // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire  [21:0] rsp_xbar_demux_004_src1_channel;                                                                     // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src1_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [93:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire  [21:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_005_src1_endofpacket;                                                                 // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src1_valid;                                                                       // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src1_startofpacket;                                                               // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [93:0] rsp_xbar_demux_005_src1_data;                                                                        // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire  [21:0] rsp_xbar_demux_005_src1_channel;                                                                     // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src1_ready;                                                                       // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [93:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	wire  [21:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_006_src1_endofpacket;                                                                 // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src1_valid;                                                                       // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src1_startofpacket;                                                               // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [93:0] rsp_xbar_demux_006_src1_data;                                                                        // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	wire  [21:0] rsp_xbar_demux_006_src1_channel;                                                                     // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src1_ready;                                                                       // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [93:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire  [21:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                       // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_007_src1_endofpacket;                                                                 // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src1_valid;                                                                       // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src1_startofpacket;                                                               // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [93:0] rsp_xbar_demux_007_src1_data;                                                                        // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire  [21:0] rsp_xbar_demux_007_src1_channel;                                                                     // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src1_ready;                                                                       // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [93:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire  [21:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                       // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_008_src1_endofpacket;                                                                 // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src1_valid;                                                                       // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src1_startofpacket;                                                               // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [93:0] rsp_xbar_demux_008_src1_data;                                                                        // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	wire  [21:0] rsp_xbar_demux_008_src1_channel;                                                                     // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src1_ready;                                                                       // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [93:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire  [21:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                       // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_009_src1_endofpacket;                                                                 // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src1_valid;                                                                       // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src1_startofpacket;                                                               // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [93:0] rsp_xbar_demux_009_src1_data;                                                                        // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	wire  [21:0] rsp_xbar_demux_009_src1_channel;                                                                     // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src1_ready;                                                                       // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [93:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire  [21:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                       // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_010_src1_endofpacket;                                                                 // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src1_valid;                                                                       // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src1_startofpacket;                                                               // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [93:0] rsp_xbar_demux_010_src1_data;                                                                        // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	wire  [21:0] rsp_xbar_demux_010_src1_channel;                                                                     // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src1_ready;                                                                       // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                                 // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                       // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                               // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [93:0] rsp_xbar_demux_011_src0_data;                                                                        // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire  [21:0] rsp_xbar_demux_011_src0_channel;                                                                     // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                       // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_011_src1_endofpacket;                                                                 // rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src1_valid;                                                                       // rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src1_startofpacket;                                                               // rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [93:0] rsp_xbar_demux_011_src1_data;                                                                        // rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_001:sink11_data
	wire  [21:0] rsp_xbar_demux_011_src1_channel;                                                                     // rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src1_ready;                                                                       // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src1_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                                 // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                       // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                               // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [93:0] rsp_xbar_demux_012_src0_data;                                                                        // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire  [21:0] rsp_xbar_demux_012_src0_channel;                                                                     // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                       // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_012_src1_endofpacket;                                                                 // rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src1_valid;                                                                       // rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src1_startofpacket;                                                               // rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [93:0] rsp_xbar_demux_012_src1_data;                                                                        // rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_001:sink12_data
	wire  [21:0] rsp_xbar_demux_012_src1_channel;                                                                     // rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src1_ready;                                                                       // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src1_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                                 // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                       // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                               // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [93:0] rsp_xbar_demux_013_src0_data;                                                                        // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire  [21:0] rsp_xbar_demux_013_src0_channel;                                                                     // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                       // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         rsp_xbar_demux_013_src1_endofpacket;                                                                 // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src1_valid;                                                                       // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src1_startofpacket;                                                               // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [93:0] rsp_xbar_demux_013_src1_data;                                                                        // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink13_data
	wire  [21:0] rsp_xbar_demux_013_src1_channel;                                                                     // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src1_ready;                                                                       // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src1_ready
	wire         rsp_xbar_demux_014_src0_endofpacket;                                                                 // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire         rsp_xbar_demux_014_src0_valid;                                                                       // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire         rsp_xbar_demux_014_src0_startofpacket;                                                               // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [93:0] rsp_xbar_demux_014_src0_data;                                                                        // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire  [21:0] rsp_xbar_demux_014_src0_channel;                                                                     // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire         rsp_xbar_demux_014_src0_ready;                                                                       // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire         rsp_xbar_demux_014_src1_endofpacket;                                                                 // rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire         rsp_xbar_demux_014_src1_valid;                                                                       // rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_001:sink14_valid
	wire         rsp_xbar_demux_014_src1_startofpacket;                                                               // rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [93:0] rsp_xbar_demux_014_src1_data;                                                                        // rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_001:sink14_data
	wire  [21:0] rsp_xbar_demux_014_src1_channel;                                                                     // rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_001:sink14_channel
	wire         rsp_xbar_demux_014_src1_ready;                                                                       // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src1_ready
	wire         rsp_xbar_demux_015_src0_endofpacket;                                                                 // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire         rsp_xbar_demux_015_src0_valid;                                                                       // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux:sink15_valid
	wire         rsp_xbar_demux_015_src0_startofpacket;                                                               // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [93:0] rsp_xbar_demux_015_src0_data;                                                                        // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux:sink15_data
	wire  [21:0] rsp_xbar_demux_015_src0_channel;                                                                     // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux:sink15_channel
	wire         rsp_xbar_demux_015_src0_ready;                                                                       // rsp_xbar_mux:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire         rsp_xbar_demux_015_src1_endofpacket;                                                                 // rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire         rsp_xbar_demux_015_src1_valid;                                                                       // rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_001:sink15_valid
	wire         rsp_xbar_demux_015_src1_startofpacket;                                                               // rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [93:0] rsp_xbar_demux_015_src1_data;                                                                        // rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_001:sink15_data
	wire  [21:0] rsp_xbar_demux_015_src1_channel;                                                                     // rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_001:sink15_channel
	wire         rsp_xbar_demux_015_src1_ready;                                                                       // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src1_ready
	wire         rsp_xbar_demux_016_src0_endofpacket;                                                                 // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	wire         rsp_xbar_demux_016_src0_valid;                                                                       // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	wire         rsp_xbar_demux_016_src0_startofpacket;                                                               // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	wire  [93:0] rsp_xbar_demux_016_src0_data;                                                                        // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	wire  [21:0] rsp_xbar_demux_016_src0_channel;                                                                     // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	wire         rsp_xbar_demux_016_src0_ready;                                                                       // rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire         rsp_xbar_demux_016_src1_endofpacket;                                                                 // rsp_xbar_demux_016:src1_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire         rsp_xbar_demux_016_src1_valid;                                                                       // rsp_xbar_demux_016:src1_valid -> rsp_xbar_mux_001:sink16_valid
	wire         rsp_xbar_demux_016_src1_startofpacket;                                                               // rsp_xbar_demux_016:src1_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [93:0] rsp_xbar_demux_016_src1_data;                                                                        // rsp_xbar_demux_016:src1_data -> rsp_xbar_mux_001:sink16_data
	wire  [21:0] rsp_xbar_demux_016_src1_channel;                                                                     // rsp_xbar_demux_016:src1_channel -> rsp_xbar_mux_001:sink16_channel
	wire         rsp_xbar_demux_016_src1_ready;                                                                       // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src1_ready
	wire         rsp_xbar_demux_017_src0_endofpacket;                                                                 // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	wire         rsp_xbar_demux_017_src0_valid;                                                                       // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	wire         rsp_xbar_demux_017_src0_startofpacket;                                                               // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	wire  [93:0] rsp_xbar_demux_017_src0_data;                                                                        // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	wire  [21:0] rsp_xbar_demux_017_src0_channel;                                                                     // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	wire         rsp_xbar_demux_017_src0_ready;                                                                       // rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire         rsp_xbar_demux_017_src1_endofpacket;                                                                 // rsp_xbar_demux_017:src1_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire         rsp_xbar_demux_017_src1_valid;                                                                       // rsp_xbar_demux_017:src1_valid -> rsp_xbar_mux_001:sink17_valid
	wire         rsp_xbar_demux_017_src1_startofpacket;                                                               // rsp_xbar_demux_017:src1_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [93:0] rsp_xbar_demux_017_src1_data;                                                                        // rsp_xbar_demux_017:src1_data -> rsp_xbar_mux_001:sink17_data
	wire  [21:0] rsp_xbar_demux_017_src1_channel;                                                                     // rsp_xbar_demux_017:src1_channel -> rsp_xbar_mux_001:sink17_channel
	wire         rsp_xbar_demux_017_src1_ready;                                                                       // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src1_ready
	wire         rsp_xbar_demux_018_src0_endofpacket;                                                                 // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	wire         rsp_xbar_demux_018_src0_valid;                                                                       // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux:sink18_valid
	wire         rsp_xbar_demux_018_src0_startofpacket;                                                               // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	wire  [93:0] rsp_xbar_demux_018_src0_data;                                                                        // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux:sink18_data
	wire  [21:0] rsp_xbar_demux_018_src0_channel;                                                                     // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux:sink18_channel
	wire         rsp_xbar_demux_018_src0_ready;                                                                       // rsp_xbar_mux:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire         rsp_xbar_demux_018_src1_endofpacket;                                                                 // rsp_xbar_demux_018:src1_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire         rsp_xbar_demux_018_src1_valid;                                                                       // rsp_xbar_demux_018:src1_valid -> rsp_xbar_mux_001:sink18_valid
	wire         rsp_xbar_demux_018_src1_startofpacket;                                                               // rsp_xbar_demux_018:src1_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [93:0] rsp_xbar_demux_018_src1_data;                                                                        // rsp_xbar_demux_018:src1_data -> rsp_xbar_mux_001:sink18_data
	wire  [21:0] rsp_xbar_demux_018_src1_channel;                                                                     // rsp_xbar_demux_018:src1_channel -> rsp_xbar_mux_001:sink18_channel
	wire         rsp_xbar_demux_018_src1_ready;                                                                       // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src1_ready
	wire         rsp_xbar_demux_019_src0_endofpacket;                                                                 // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux:sink19_endofpacket
	wire         rsp_xbar_demux_019_src0_valid;                                                                       // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux:sink19_valid
	wire         rsp_xbar_demux_019_src0_startofpacket;                                                               // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux:sink19_startofpacket
	wire  [93:0] rsp_xbar_demux_019_src0_data;                                                                        // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux:sink19_data
	wire  [21:0] rsp_xbar_demux_019_src0_channel;                                                                     // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux:sink19_channel
	wire         rsp_xbar_demux_019_src0_ready;                                                                       // rsp_xbar_mux:sink19_ready -> rsp_xbar_demux_019:src0_ready
	wire         rsp_xbar_demux_019_src1_endofpacket;                                                                 // rsp_xbar_demux_019:src1_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	wire         rsp_xbar_demux_019_src1_valid;                                                                       // rsp_xbar_demux_019:src1_valid -> rsp_xbar_mux_001:sink19_valid
	wire         rsp_xbar_demux_019_src1_startofpacket;                                                               // rsp_xbar_demux_019:src1_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	wire  [93:0] rsp_xbar_demux_019_src1_data;                                                                        // rsp_xbar_demux_019:src1_data -> rsp_xbar_mux_001:sink19_data
	wire  [21:0] rsp_xbar_demux_019_src1_channel;                                                                     // rsp_xbar_demux_019:src1_channel -> rsp_xbar_mux_001:sink19_channel
	wire         rsp_xbar_demux_019_src1_ready;                                                                       // rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src1_ready
	wire         rsp_xbar_demux_020_src0_endofpacket;                                                                 // rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux:sink20_endofpacket
	wire         rsp_xbar_demux_020_src0_valid;                                                                       // rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux:sink20_valid
	wire         rsp_xbar_demux_020_src0_startofpacket;                                                               // rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux:sink20_startofpacket
	wire  [93:0] rsp_xbar_demux_020_src0_data;                                                                        // rsp_xbar_demux_020:src0_data -> rsp_xbar_mux:sink20_data
	wire  [21:0] rsp_xbar_demux_020_src0_channel;                                                                     // rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux:sink20_channel
	wire         rsp_xbar_demux_020_src0_ready;                                                                       // rsp_xbar_mux:sink20_ready -> rsp_xbar_demux_020:src0_ready
	wire         rsp_xbar_demux_020_src1_endofpacket;                                                                 // rsp_xbar_demux_020:src1_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	wire         rsp_xbar_demux_020_src1_valid;                                                                       // rsp_xbar_demux_020:src1_valid -> rsp_xbar_mux_001:sink20_valid
	wire         rsp_xbar_demux_020_src1_startofpacket;                                                               // rsp_xbar_demux_020:src1_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	wire  [93:0] rsp_xbar_demux_020_src1_data;                                                                        // rsp_xbar_demux_020:src1_data -> rsp_xbar_mux_001:sink20_data
	wire  [21:0] rsp_xbar_demux_020_src1_channel;                                                                     // rsp_xbar_demux_020:src1_channel -> rsp_xbar_mux_001:sink20_channel
	wire         rsp_xbar_demux_020_src1_ready;                                                                       // rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src1_ready
	wire         rsp_xbar_demux_021_src0_endofpacket;                                                                 // rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux:sink21_endofpacket
	wire         rsp_xbar_demux_021_src0_valid;                                                                       // rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux:sink21_valid
	wire         rsp_xbar_demux_021_src0_startofpacket;                                                               // rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux:sink21_startofpacket
	wire  [93:0] rsp_xbar_demux_021_src0_data;                                                                        // rsp_xbar_demux_021:src0_data -> rsp_xbar_mux:sink21_data
	wire  [21:0] rsp_xbar_demux_021_src0_channel;                                                                     // rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux:sink21_channel
	wire         rsp_xbar_demux_021_src0_ready;                                                                       // rsp_xbar_mux:sink21_ready -> rsp_xbar_demux_021:src0_ready
	wire         rsp_xbar_demux_021_src1_endofpacket;                                                                 // rsp_xbar_demux_021:src1_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	wire         rsp_xbar_demux_021_src1_valid;                                                                       // rsp_xbar_demux_021:src1_valid -> rsp_xbar_mux_001:sink21_valid
	wire         rsp_xbar_demux_021_src1_startofpacket;                                                               // rsp_xbar_demux_021:src1_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	wire  [93:0] rsp_xbar_demux_021_src1_data;                                                                        // rsp_xbar_demux_021:src1_data -> rsp_xbar_mux_001:sink21_data
	wire  [21:0] rsp_xbar_demux_021_src1_channel;                                                                     // rsp_xbar_demux_021:src1_channel -> rsp_xbar_mux_001:sink21_channel
	wire         rsp_xbar_demux_021_src1_ready;                                                                       // rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src1_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [93:0] addr_router_src_data;                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire  [21:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [21:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [93:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire  [21:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [93:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [21:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [93:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [21:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [93:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [21:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                             // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                          // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [93:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [21:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_mux_003_src_endofpacket;                                                                    // cmd_xbar_mux_003:src_endofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_003_src_valid;                                                                          // cmd_xbar_mux_003:src_valid -> switch_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_003_src_startofpacket;                                                                  // cmd_xbar_mux_003:src_startofpacket -> switch_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_003_src_data;                                                                           // cmd_xbar_mux_003:src_data -> switch_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_003_src_channel;                                                                        // cmd_xbar_mux_003:src_channel -> switch_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_003_src_ready;                                                                          // switch_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [93:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [21:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_mux_004_src_endofpacket;                                                                    // cmd_xbar_mux_004:src_endofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_004_src_valid;                                                                          // cmd_xbar_mux_004:src_valid -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_004_src_startofpacket;                                                                  // cmd_xbar_mux_004:src_startofpacket -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_004_src_data;                                                                           // cmd_xbar_mux_004:src_data -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_004_src_channel;                                                                        // cmd_xbar_mux_004:src_channel -> ledr_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_004_src_ready;                                                                          // ledr_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [93:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [21:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_mux_005_src_endofpacket;                                                                    // cmd_xbar_mux_005:src_endofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_005_src_valid;                                                                          // cmd_xbar_mux_005:src_valid -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_005_src_startofpacket;                                                                  // cmd_xbar_mux_005:src_startofpacket -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_005_src_data;                                                                           // cmd_xbar_mux_005:src_data -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_005_src_channel;                                                                        // cmd_xbar_mux_005:src_channel -> hex0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_005_src_ready;                                                                          // hex0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [93:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [21:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_006_src_endofpacket;                                                                    // cmd_xbar_mux_006:src_endofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_006_src_valid;                                                                          // cmd_xbar_mux_006:src_valid -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_006_src_startofpacket;                                                                  // cmd_xbar_mux_006:src_startofpacket -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_006_src_data;                                                                           // cmd_xbar_mux_006:src_data -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_006_src_channel;                                                                        // cmd_xbar_mux_006:src_channel -> hex1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_006_src_ready;                                                                          // hex1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	wire         id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [93:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [21:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_mux_007_src_endofpacket;                                                                    // cmd_xbar_mux_007:src_endofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_007_src_valid;                                                                          // cmd_xbar_mux_007:src_valid -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_007_src_startofpacket;                                                                  // cmd_xbar_mux_007:src_startofpacket -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_007_src_data;                                                                           // cmd_xbar_mux_007:src_data -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_007_src_channel;                                                                        // cmd_xbar_mux_007:src_channel -> hex2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_007_src_ready;                                                                          // hex2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire         id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [93:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [21:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_mux_008_src_endofpacket;                                                                    // cmd_xbar_mux_008:src_endofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_008_src_valid;                                                                          // cmd_xbar_mux_008:src_valid -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_008_src_startofpacket;                                                                  // cmd_xbar_mux_008:src_startofpacket -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_008_src_data;                                                                           // cmd_xbar_mux_008:src_data -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_008_src_channel;                                                                        // cmd_xbar_mux_008:src_channel -> hex3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_008_src_ready;                                                                          // hex3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire         id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [93:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [21:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_mux_009_src_endofpacket;                                                                    // cmd_xbar_mux_009:src_endofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_009_src_valid;                                                                          // cmd_xbar_mux_009:src_valid -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_009_src_startofpacket;                                                                  // cmd_xbar_mux_009:src_startofpacket -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_009_src_data;                                                                           // cmd_xbar_mux_009:src_data -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_009_src_channel;                                                                        // cmd_xbar_mux_009:src_channel -> hex4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_009_src_ready;                                                                          // hex4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire         id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [93:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [21:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_mux_010_src_endofpacket;                                                                    // cmd_xbar_mux_010:src_endofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_010_src_valid;                                                                          // cmd_xbar_mux_010:src_valid -> hex5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_010_src_startofpacket;                                                                  // cmd_xbar_mux_010:src_startofpacket -> hex5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_010_src_data;                                                                           // cmd_xbar_mux_010:src_data -> hex5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_010_src_channel;                                                                        // cmd_xbar_mux_010:src_channel -> hex5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_010_src_ready;                                                                          // hex5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire         id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                             // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [93:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [21:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                             // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_mux_011_src_endofpacket;                                                                    // cmd_xbar_mux_011:src_endofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_011_src_valid;                                                                          // cmd_xbar_mux_011:src_valid -> hex6_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_011_src_startofpacket;                                                                  // cmd_xbar_mux_011:src_startofpacket -> hex6_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_011_src_data;                                                                           // cmd_xbar_mux_011:src_data -> hex6_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_011_src_channel;                                                                        // cmd_xbar_mux_011:src_channel -> hex6_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_011_src_ready;                                                                          // hex6_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	wire         id_router_011_src_endofpacket;                                                                       // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                             // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                     // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [93:0] id_router_011_src_data;                                                                              // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [21:0] id_router_011_src_channel;                                                                           // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                             // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_mux_012_src_endofpacket;                                                                    // cmd_xbar_mux_012:src_endofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_012_src_valid;                                                                          // cmd_xbar_mux_012:src_valid -> hex7_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_012_src_startofpacket;                                                                  // cmd_xbar_mux_012:src_startofpacket -> hex7_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_012_src_data;                                                                           // cmd_xbar_mux_012:src_data -> hex7_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_012_src_channel;                                                                        // cmd_xbar_mux_012:src_channel -> hex7_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_012_src_ready;                                                                          // hex7_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	wire         id_router_012_src_endofpacket;                                                                       // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                             // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                     // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [93:0] id_router_012_src_data;                                                                              // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [21:0] id_router_012_src_channel;                                                                           // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                             // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_mux_013_src_endofpacket;                                                                    // cmd_xbar_mux_013:src_endofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_013_src_valid;                                                                          // cmd_xbar_mux_013:src_valid -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_013_src_startofpacket;                                                                  // cmd_xbar_mux_013:src_startofpacket -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_013_src_data;                                                                           // cmd_xbar_mux_013:src_data -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_013_src_channel;                                                                        // cmd_xbar_mux_013:src_channel -> ledg_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_013_src_ready;                                                                          // ledg_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire         id_router_013_src_endofpacket;                                                                       // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                             // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                     // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [93:0] id_router_013_src_data;                                                                              // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [21:0] id_router_013_src_channel;                                                                           // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                             // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire         cmd_xbar_mux_014_src_endofpacket;                                                                    // cmd_xbar_mux_014:src_endofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_014_src_valid;                                                                          // cmd_xbar_mux_014:src_valid -> key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_014_src_startofpacket;                                                                  // cmd_xbar_mux_014:src_startofpacket -> key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_014_src_data;                                                                           // cmd_xbar_mux_014:src_data -> key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_014_src_channel;                                                                        // cmd_xbar_mux_014:src_channel -> key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_014_src_ready;                                                                          // key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	wire         id_router_014_src_endofpacket;                                                                       // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire         id_router_014_src_valid;                                                                             // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire         id_router_014_src_startofpacket;                                                                     // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [93:0] id_router_014_src_data;                                                                              // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire  [21:0] id_router_014_src_channel;                                                                           // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire         id_router_014_src_ready;                                                                             // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire         cmd_xbar_mux_015_src_endofpacket;                                                                    // cmd_xbar_mux_015:src_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_015_src_valid;                                                                          // cmd_xbar_mux_015:src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_015_src_startofpacket;                                                                  // cmd_xbar_mux_015:src_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_015_src_data;                                                                           // cmd_xbar_mux_015:src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_015_src_channel;                                                                        // cmd_xbar_mux_015:src_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_015_src_ready;                                                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	wire         id_router_015_src_endofpacket;                                                                       // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire         id_router_015_src_valid;                                                                             // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire         id_router_015_src_startofpacket;                                                                     // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [93:0] id_router_015_src_data;                                                                              // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire  [21:0] id_router_015_src_channel;                                                                           // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire         id_router_015_src_ready;                                                                             // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire         cmd_xbar_mux_016_src_endofpacket;                                                                    // cmd_xbar_mux_016:src_endofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_016_src_valid;                                                                          // cmd_xbar_mux_016:src_valid -> lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_016_src_startofpacket;                                                                  // cmd_xbar_mux_016:src_startofpacket -> lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_016_src_data;                                                                           // cmd_xbar_mux_016:src_data -> lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_016_src_channel;                                                                        // cmd_xbar_mux_016:src_channel -> lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_016_src_ready;                                                                          // lcd_d_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_016:src_ready
	wire         id_router_016_src_endofpacket;                                                                       // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire         id_router_016_src_valid;                                                                             // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire         id_router_016_src_startofpacket;                                                                     // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [93:0] id_router_016_src_data;                                                                              // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire  [21:0] id_router_016_src_channel;                                                                           // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire         id_router_016_src_ready;                                                                             // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire         cmd_xbar_mux_017_src_endofpacket;                                                                    // cmd_xbar_mux_017:src_endofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_017_src_valid;                                                                          // cmd_xbar_mux_017:src_valid -> lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_017_src_startofpacket;                                                                  // cmd_xbar_mux_017:src_startofpacket -> lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_017_src_data;                                                                           // cmd_xbar_mux_017:src_data -> lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_017_src_channel;                                                                        // cmd_xbar_mux_017:src_channel -> lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_017_src_ready;                                                                          // lcd_on_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_017:src_ready
	wire         id_router_017_src_endofpacket;                                                                       // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire         id_router_017_src_valid;                                                                             // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire         id_router_017_src_startofpacket;                                                                     // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [93:0] id_router_017_src_data;                                                                              // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire  [21:0] id_router_017_src_channel;                                                                           // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire         id_router_017_src_ready;                                                                             // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire         cmd_xbar_mux_018_src_endofpacket;                                                                    // cmd_xbar_mux_018:src_endofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_018_src_valid;                                                                          // cmd_xbar_mux_018:src_valid -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_018_src_startofpacket;                                                                  // cmd_xbar_mux_018:src_startofpacket -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_018_src_data;                                                                           // cmd_xbar_mux_018:src_data -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_018_src_channel;                                                                        // cmd_xbar_mux_018:src_channel -> lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_018_src_ready;                                                                          // lcd_blon_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_018:src_ready
	wire         id_router_018_src_endofpacket;                                                                       // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire         id_router_018_src_valid;                                                                             // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire         id_router_018_src_startofpacket;                                                                     // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [93:0] id_router_018_src_data;                                                                              // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire  [21:0] id_router_018_src_channel;                                                                           // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire         id_router_018_src_ready;                                                                             // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire         cmd_xbar_mux_019_src_endofpacket;                                                                    // cmd_xbar_mux_019:src_endofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_019_src_valid;                                                                          // cmd_xbar_mux_019:src_valid -> lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_019_src_startofpacket;                                                                  // cmd_xbar_mux_019:src_startofpacket -> lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_019_src_data;                                                                           // cmd_xbar_mux_019:src_data -> lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_019_src_channel;                                                                        // cmd_xbar_mux_019:src_channel -> lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_019_src_ready;                                                                          // lcd_en_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_019:src_ready
	wire         id_router_019_src_endofpacket;                                                                       // id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire         id_router_019_src_valid;                                                                             // id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	wire         id_router_019_src_startofpacket;                                                                     // id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire  [93:0] id_router_019_src_data;                                                                              // id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	wire  [21:0] id_router_019_src_channel;                                                                           // id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	wire         id_router_019_src_ready;                                                                             // rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	wire         cmd_xbar_mux_020_src_endofpacket;                                                                    // cmd_xbar_mux_020:src_endofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_020_src_valid;                                                                          // cmd_xbar_mux_020:src_valid -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_020_src_startofpacket;                                                                  // cmd_xbar_mux_020:src_startofpacket -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_020_src_data;                                                                           // cmd_xbar_mux_020:src_data -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_020_src_channel;                                                                        // cmd_xbar_mux_020:src_channel -> lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_020_src_ready;                                                                          // lcd_rw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_020:src_ready
	wire         id_router_020_src_endofpacket;                                                                       // id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire         id_router_020_src_valid;                                                                             // id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	wire         id_router_020_src_startofpacket;                                                                     // id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [93:0] id_router_020_src_data;                                                                              // id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	wire  [21:0] id_router_020_src_channel;                                                                           // id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	wire         id_router_020_src_ready;                                                                             // rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	wire         cmd_xbar_mux_021_src_endofpacket;                                                                    // cmd_xbar_mux_021:src_endofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_021_src_valid;                                                                          // cmd_xbar_mux_021:src_valid -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_021_src_startofpacket;                                                                  // cmd_xbar_mux_021:src_startofpacket -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [93:0] cmd_xbar_mux_021_src_data;                                                                           // cmd_xbar_mux_021:src_data -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [21:0] cmd_xbar_mux_021_src_channel;                                                                        // cmd_xbar_mux_021:src_channel -> lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_021_src_ready;                                                                          // lcd_rs_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_021:src_ready
	wire         id_router_021_src_endofpacket;                                                                       // id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	wire         id_router_021_src_valid;                                                                             // id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	wire         id_router_021_src_startofpacket;                                                                     // id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	wire  [93:0] id_router_021_src_data;                                                                              // id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	wire  [21:0] id_router_021_src_channel;                                                                           // id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	wire         id_router_021_src_ready;                                                                             // rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	wire         irq_mapper_receiver0_irq;                                                                            // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                            // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	nios_sys_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (clk_clk),                                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	nios_sys_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                                       //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                             //       .reset_req
	);

	nios_sys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_sys_switch switch (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (switch_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (switch_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switch_external_connection_export)                  // external_connection.export
	);

	nios_sys_ledr ledr (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledr_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex0 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex0_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex0_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex0_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex0_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex0_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex0_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex1 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex1_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex2 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex2_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex3 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex3_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex3_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex3_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex3_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex3_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex3_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex4 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex4_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex4_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex4_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex4_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex4_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex4_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex5 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex5_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex5_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex5_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex5_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex5_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex5_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex6 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex6_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex6_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex6_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex6_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex6_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex6_external_connection_export)                    // external_connection.export
	);

	nios_sys_hex0 hex7 (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (hex7_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hex7_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hex7_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hex7_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hex7_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex7_external_connection_export)                    // external_connection.export
	);

	nios_sys_ledg ledg (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (ledg_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~ledg_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (ledg_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (ledg_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (ledg_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (ledg_external_connection_export)                    // external_connection.export
	);

	nios_sys_key key (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (key_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (key_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (key_external_connection_export)                  // external_connection.export
	);

	nios_sys_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                              //   irq.irq
	);

	nios_sys_lcd_d lcd_d (
		.clk        (clk_clk),                                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (lcd_d_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_d_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_d_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_d_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_d_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_d_external_connection_export)                    // external_connection.export
	);

	nios_sys_lcd_on lcd_on (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_on_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_on_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_on_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_on_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_on_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_on_external_connection_export)                    // external_connection.export
	);

	nios_sys_lcd_on lcd_blon (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (lcd_blon_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_blon_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_blon_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_blon_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_blon_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_blon_external_connection_export)                    // external_connection.export
	);

	nios_sys_lcd_on lcd_en (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_en_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_en_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_en_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_en_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_en_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_en_external_connection_export)                    // external_connection.export
	);

	nios_sys_lcd_on lcd_rw (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_rw_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_rw_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_rw_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_rw_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_rw_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_rw_external_connection_export)                    // external_connection.export
	);

	nios_sys_lcd_on lcd_rs (
		.clk        (clk_clk),                                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_rs_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_rs_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_rs_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_rs_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_rs_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (lcd_rs_external_connection_export)                    // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (17),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (17),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (clk_clk),                                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_readdatavalid         (),                                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (17),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (17),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                      (clk_clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (13),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (clk_clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) switch_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (switch_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (switch_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                     //              (terminated)
		.av_read                  (),                                                                     //              (terminated)
		.av_writedata             (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_chipselect            (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledr_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex0_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex1_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex2_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex3_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex4_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex5_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex6_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex6_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex6_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex6_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex6_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex6_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex6_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex6_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex6_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex6_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hex7_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (hex7_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (hex7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (hex7_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (hex7_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (hex7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (hex7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (hex7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (hex7_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (hex7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (hex7_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (hex7_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (hex7_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (hex7_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (hex7_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ledg_s1_translator (
		.clk                      (clk_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ledg_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ledg_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ledg_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ledg_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (ledg_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                   //              (terminated)
		.av_begintransfer         (),                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                   //              (terminated)
		.av_burstcount            (),                                                                   //              (terminated)
		.av_byteenable            (),                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                               //              (terminated)
		.av_writebyteenable       (),                                                                   //              (terminated)
		.av_lock                  (),                                                                   //              (terminated)
		.av_clken                 (),                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                               //              (terminated)
		.av_debugaccess           (),                                                                   //              (terminated)
		.av_outputenable          (),                                                                   //              (terminated)
		.uav_response             (),                                                                   //              (terminated)
		.av_response              (2'b00),                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) key_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                  //              (terminated)
		.av_read                  (),                                                                  //              (terminated)
		.av_writedata             (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_byteenable            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.av_chipselect            (),                                                                  //              (terminated)
		.av_clken                 (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_d_s1_translator (
		.clk                      (clk_clk),                                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_d_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_d_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_d_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_d_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_d_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_on_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_on_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_on_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_on_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_on_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_on_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_blon_s1_translator (
		.clk                      (clk_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_blon_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_blon_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_blon_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_blon_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_blon_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_en_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_en_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_en_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_en_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_en_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_en_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_rw_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_rw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_rw_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_rw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_rw_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_rw_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (17),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_rs_s1_translator (
		.clk                      (clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_rs_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_rs_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_rs_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_rs_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_rs_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                     //              (terminated)
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_burstcount            (),                                                                     //              (terminated)
		.av_byteenable            (),                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_lock                  (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_debugaccess           (),                                                                     //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.PKT_BURST_TYPE_H          (69),
		.PKT_BURST_TYPE_L          (68),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_TRANS_EXCLUSIVE       (58),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (71),
		.PKT_DATA_SIDEBAND_L       (71),
		.PKT_QOS_H                 (73),
		.PKT_QOS_L                 (73),
		.PKT_ADDR_SIDEBAND_H       (70),
		.PKT_ADDR_SIDEBAND_L       (70),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (22),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                       //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                      //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (72),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.PKT_BURST_TYPE_H          (69),
		.PKT_BURST_TYPE_L          (68),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_TRANS_EXCLUSIVE       (58),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (71),
		.PKT_DATA_SIDEBAND_L       (71),
		.PKT_QOS_H                 (73),
		.PKT_QOS_L                 (73),
		.PKT_ADDR_SIDEBAND_H       (70),
		.PKT_ADDR_SIDEBAND_L       (70),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (22),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                            //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                           //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                       //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) switch_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (switch_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (switch_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (switch_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (switch_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (switch_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (switch_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (switch_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (switch_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (switch_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                   //                .channel
		.rf_sink_ready           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (switch_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (switch_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                 //                .channel
		.rf_sink_ready           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_006_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_006_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_006_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_006_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_006_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_006_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex6_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex6_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex6_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex6_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex6_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex6_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex6_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex6_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_011_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_011_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_011_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_011_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_011_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_011_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) hex7_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (hex7_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hex7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hex7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hex7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hex7_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hex7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hex7_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hex7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hex7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hex7_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hex7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hex7_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hex7_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hex7_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hex7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_012_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_012_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_012_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_012_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_012_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_012_src_channel),                                                 //                .channel
		.rf_sink_ready           (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hex7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hex7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hex7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                 //                .channel
		.rf_sink_ready           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_014_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_014_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_014_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_014_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_014_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_014_src_channel),                                                //                .channel
		.rf_sink_ready           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_015_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_015_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_015_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_015_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_015_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_015_src_channel),                                                    //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_d_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_d_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_016_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_016_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_016_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_016_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_016_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_016_src_channel),                                                  //                .channel
		.rf_sink_ready           (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_d_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_d_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_on_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_on_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_017_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_017_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_017_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_017_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_017_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_017_src_channel),                                                   //                .channel
		.rf_sink_ready           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_on_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_on_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_blon_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_blon_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_018_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_018_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_018_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_018_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_018_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_018_src_channel),                                                     //                .channel
		.rf_sink_ready           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_en_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_en_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_019_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_019_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_019_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_019_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_019_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_019_src_channel),                                                   //                .channel
		.rf_sink_ready           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_rw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_020_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_020_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_020_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_020_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_020_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_020_src_channel),                                                   //                .channel
		.rf_sink_ready           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (72),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (52),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (53),
		.PKT_TRANS_POSTED          (54),
		.PKT_TRANS_WRITE           (55),
		.PKT_TRANS_READ            (56),
		.PKT_TRANS_LOCK            (57),
		.PKT_SRC_ID_H              (78),
		.PKT_SRC_ID_L              (74),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (79),
		.PKT_BURSTWRAP_H           (64),
		.PKT_BURSTWRAP_L           (62),
		.PKT_BYTE_CNT_H            (61),
		.PKT_BYTE_CNT_L            (59),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (67),
		.PKT_BURST_SIZE_L          (65),
		.ST_CHANNEL_W              (22),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_rs_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_021_src_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_021_src_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_021_src_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_021_src_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_021_src_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_021_src_channel),                                                   //                .channel
		.rf_sink_ready           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	nios_sys_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_sys_addr_router addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios_sys_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_sys_id_router id_router_001 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                             //          .endofpacket
	);

	nios_sys_id_router id_router_002 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                        //       src.ready
		.src_valid          (id_router_002_src_valid),                                                        //          .valid
		.src_data           (id_router_002_src_data),                                                         //          .data
		.src_channel        (id_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	nios_sys_id_router id_router_003 (
		.sink_ready         (switch_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (switch_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (switch_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (switch_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (switch_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                              //       src.ready
		.src_valid          (id_router_003_src_valid),                                              //          .valid
		.src_data           (id_router_003_src_data),                                               //          .data
		.src_channel        (id_router_003_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router id_router_004 (
		.sink_ready         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                            //       src.ready
		.src_valid          (id_router_004_src_valid),                                            //          .valid
		.src_data           (id_router_004_src_data),                                             //          .data
		.src_channel        (id_router_004_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_005 (
		.sink_ready         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                            //       src.ready
		.src_valid          (id_router_005_src_valid),                                            //          .valid
		.src_data           (id_router_005_src_data),                                             //          .data
		.src_channel        (id_router_005_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_006 (
		.sink_ready         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                            //       src.ready
		.src_valid          (id_router_006_src_valid),                                            //          .valid
		.src_data           (id_router_006_src_data),                                             //          .data
		.src_channel        (id_router_006_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_007 (
		.sink_ready         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                            //       src.ready
		.src_valid          (id_router_007_src_valid),                                            //          .valid
		.src_data           (id_router_007_src_data),                                             //          .data
		.src_channel        (id_router_007_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_008 (
		.sink_ready         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                            //       src.ready
		.src_valid          (id_router_008_src_valid),                                            //          .valid
		.src_data           (id_router_008_src_data),                                             //          .data
		.src_channel        (id_router_008_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_009 (
		.sink_ready         (hex4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                            //          .valid
		.src_data           (id_router_009_src_data),                                             //          .data
		.src_channel        (id_router_009_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_010 (
		.sink_ready         (hex5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                            //       src.ready
		.src_valid          (id_router_010_src_valid),                                            //          .valid
		.src_data           (id_router_010_src_data),                                             //          .data
		.src_channel        (id_router_010_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_011 (
		.sink_ready         (hex6_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex6_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex6_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                            //       src.ready
		.src_valid          (id_router_011_src_valid),                                            //          .valid
		.src_data           (id_router_011_src_data),                                             //          .data
		.src_channel        (id_router_011_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_012 (
		.sink_ready         (hex7_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hex7_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hex7_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hex7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hex7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                            //       src.ready
		.src_valid          (id_router_012_src_valid),                                            //          .valid
		.src_data           (id_router_012_src_data),                                             //          .data
		.src_channel        (id_router_012_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_013 (
		.sink_ready         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                            //       src.ready
		.src_valid          (id_router_013_src_valid),                                            //          .valid
		.src_data           (id_router_013_src_data),                                             //          .data
		.src_channel        (id_router_013_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                       //          .endofpacket
	);

	nios_sys_id_router id_router_014 (
		.sink_ready         (key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                           //       src.ready
		.src_valid          (id_router_014_src_valid),                                           //          .valid
		.src_data           (id_router_014_src_data),                                            //          .data
		.src_channel        (id_router_014_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                      //          .endofpacket
	);

	nios_sys_id_router id_router_015 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	nios_sys_id_router id_router_016 (
		.sink_ready         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_d_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                             //       src.ready
		.src_valid          (id_router_016_src_valid),                                             //          .valid
		.src_data           (id_router_016_src_data),                                              //          .data
		.src_channel        (id_router_016_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                        //          .endofpacket
	);

	nios_sys_id_router id_router_017 (
		.sink_ready         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_on_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                              //       src.ready
		.src_valid          (id_router_017_src_valid),                                              //          .valid
		.src_data           (id_router_017_src_data),                                               //          .data
		.src_channel        (id_router_017_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router id_router_018 (
		.sink_ready         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_blon_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                //       src.ready
		.src_valid          (id_router_018_src_valid),                                                //          .valid
		.src_data           (id_router_018_src_data),                                                 //          .data
		.src_channel        (id_router_018_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                           //          .endofpacket
	);

	nios_sys_id_router id_router_019 (
		.sink_ready         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                              //       src.ready
		.src_valid          (id_router_019_src_valid),                                              //          .valid
		.src_data           (id_router_019_src_data),                                               //          .data
		.src_channel        (id_router_019_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router id_router_020 (
		.sink_ready         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_rw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                              //       src.ready
		.src_valid          (id_router_020_src_valid),                                              //          .valid
		.src_data           (id_router_020_src_data),                                               //          .data
		.src_channel        (id_router_020_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                         //          .endofpacket
	);

	nios_sys_id_router id_router_021 (
		.sink_ready         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_rs_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_021_src_ready),                                              //       src.ready
		.src_valid          (id_router_021_src_valid),                                              //          .valid
		.src_data           (id_router_021_src_data),                                               //          .data
		.src_channel        (id_router_021_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_021_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_021_src_endofpacket)                                         //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	nios_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (clk_clk),                            //       clk.clk
		.reset               (rst_controller_reset_out_reset),     // clk_reset.reset
		.sink_ready          (addr_router_src_ready),              //      sink.ready
		.sink_channel        (addr_router_src_channel),            //          .channel
		.sink_data           (addr_router_src_data),               //          .data
		.sink_startofpacket  (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_src21_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //     src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //          .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //     src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //          .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //     src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket),   //          .endofpacket
		.src19_ready         (cmd_xbar_demux_001_src19_ready),         //     src19.ready
		.src19_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.src19_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.src19_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.src19_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.src19_endofpacket   (cmd_xbar_demux_001_src19_endofpacket),   //          .endofpacket
		.src20_ready         (cmd_xbar_demux_001_src20_ready),         //     src20.ready
		.src20_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.src20_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.src20_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.src20_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.src20_endofpacket   (cmd_xbar_demux_001_src20_endofpacket),   //          .endofpacket
		.src21_ready         (cmd_xbar_demux_001_src21_ready),         //     src21.ready
		.src21_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.src21_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.src21_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.src21_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.src21_endofpacket   (cmd_xbar_demux_001_src21_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src6_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src6_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src6_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src6_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src6_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src6_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src6_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src6_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src6_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src6_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src6_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src9_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src9_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src9_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src9_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src9_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src9_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src9_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src9_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src10_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src10_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src10_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src10_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src10_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src10_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src10_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_011 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_011_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_011_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src11_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src11_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src11_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src11_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src11_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src11_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src11_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src11_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_012 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src12_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src12_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src12_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src12_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src12_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src12_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src12_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src13_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src13_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src13_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src13_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src13_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src13_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src13_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src13_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_014 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_014_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_014_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_014_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_014_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_014_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_014_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src14_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src14_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src14_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src14_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src14_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src14_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src14_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src14_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_015 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src15_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src15_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src15_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src15_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src15_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src15_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src15_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src15_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_016 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_016_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_016_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_016_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_016_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_016_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_016_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src16_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src16_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src16_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src16_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src16_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src16_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src16_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src16_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src16_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src16_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src16_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_017 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_017_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_017_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_017_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_017_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_017_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_017_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src17_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src17_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src17_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src17_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src17_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src17_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src17_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src17_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src17_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src17_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src17_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_018 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_018_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_018_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_018_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_018_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_018_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_018_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src18_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src18_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src18_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src18_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src18_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src18_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src18_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src18_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src18_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src18_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src18_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_019 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_019_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_019_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_019_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_019_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_019_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_019_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src19_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src19_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src19_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src19_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src19_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src19_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src19_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src19_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src19_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src19_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src19_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src19_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_020 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_020_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_020_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_020_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_020_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_020_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_020_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src20_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src20_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src20_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src20_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src20_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src20_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src20_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src20_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src20_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src20_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src20_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src20_endofpacket)    //          .endofpacket
	);

	nios_sys_cmd_xbar_mux cmd_xbar_mux_021 (
		.clk                 (clk_clk),                                //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_021_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_021_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_021_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_021_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_021_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_021_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src21_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src21_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src21_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src21_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src21_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src21_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src21_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src21_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src21_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src21_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src21_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src21_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_011_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_014 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_014_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_015 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_016 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_016_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_016_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_017 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_017_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_017_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_018 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_018_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_018_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_019 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_019_src_ready),               //      sink.ready
		.sink_channel       (id_router_019_src_channel),             //          .channel
		.sink_data          (id_router_019_src_data),                //          .data
		.sink_startofpacket (id_router_019_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_019_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_019_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_019_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_019_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_019_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_019_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_019_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_020 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_020_src_ready),               //      sink.ready
		.sink_channel       (id_router_020_src_channel),             //          .channel
		.sink_data          (id_router_020_src_data),                //          .data
		.sink_startofpacket (id_router_020_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_020_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_020_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_020_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_020_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_020_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_020_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_020_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_020_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_demux rsp_xbar_demux_021 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_021_src_ready),               //      sink.ready
		.sink_channel       (id_router_021_src_channel),             //          .channel
		.sink_data          (id_router_021_src_data),                //          .data
		.sink_startofpacket (id_router_021_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_021_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_021_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_021_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_021_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_021_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_021_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src0_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src0_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src0_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src0_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src0_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src0_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src0_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src0_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src0_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src0_endofpacket)    //          .endofpacket
	);

	nios_sys_rsp_xbar_mux rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src1_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src1_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src1_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src1_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src1_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src1_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src1_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src1_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src1_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src1_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src1_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src1_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src1_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src1_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src1_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src1_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src1_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src1_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src1_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src1_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src1_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src1_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src1_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src1_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src1_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src1_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src1_endofpacket),   //          .endofpacket
		.sink19_ready         (rsp_xbar_demux_019_src1_ready),         //    sink19.ready
		.sink19_valid         (rsp_xbar_demux_019_src1_valid),         //          .valid
		.sink19_channel       (rsp_xbar_demux_019_src1_channel),       //          .channel
		.sink19_data          (rsp_xbar_demux_019_src1_data),          //          .data
		.sink19_startofpacket (rsp_xbar_demux_019_src1_startofpacket), //          .startofpacket
		.sink19_endofpacket   (rsp_xbar_demux_019_src1_endofpacket),   //          .endofpacket
		.sink20_ready         (rsp_xbar_demux_020_src1_ready),         //    sink20.ready
		.sink20_valid         (rsp_xbar_demux_020_src1_valid),         //          .valid
		.sink20_channel       (rsp_xbar_demux_020_src1_channel),       //          .channel
		.sink20_data          (rsp_xbar_demux_020_src1_data),          //          .data
		.sink20_startofpacket (rsp_xbar_demux_020_src1_startofpacket), //          .startofpacket
		.sink20_endofpacket   (rsp_xbar_demux_020_src1_endofpacket),   //          .endofpacket
		.sink21_ready         (rsp_xbar_demux_021_src1_ready),         //    sink21.ready
		.sink21_valid         (rsp_xbar_demux_021_src1_valid),         //          .valid
		.sink21_channel       (rsp_xbar_demux_021_src1_channel),       //          .channel
		.sink21_data          (rsp_xbar_demux_021_src1_data),          //          .data
		.sink21_startofpacket (rsp_xbar_demux_021_src1_startofpacket), //          .startofpacket
		.sink21_endofpacket   (rsp_xbar_demux_021_src1_endofpacket)    //          .endofpacket
	);

	nios_sys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
